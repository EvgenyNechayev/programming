library verilog;
use verilog.vl_types.all;
entity test_truth_table_v1 is
end test_truth_table_v1;
