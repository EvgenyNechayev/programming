library verilog;
use verilog.vl_types.all;
entity test_d_trigger is
end test_d_trigger;
