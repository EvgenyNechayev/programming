library verilog;
use verilog.vl_types.all;
entity test_simple_processor is
    generic(
        BITS            : integer := 16
    );
end test_simple_processor;
