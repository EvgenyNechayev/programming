library verilog;
use verilog.vl_types.all;
entity test_demultiplexer is
end test_demultiplexer;
