library verilog;
use verilog.vl_types.all;
entity test_par_to_ser is
    generic(
        PREAMBLE        : integer := 6
    );
end test_par_to_ser;
