
// Модуль управления сериализацией  
module control_block
	#(parameter N = 5)			// Максимально допустимое количество байт входных данных 
	(
	input  wire 	  rst_i,		// Сигнал асинхронного сброса 
	input  wire 	  clk_i,		// Синхросигнал, по которому работает модуль 
	input  wire 	  en_i,			// Сигнал валидности входных данных 
	input  wire [7:0] data_i,		// Восемь бит входных данных  
	input  wire [3:0] count_i,		// Счетчик - для проверки конца передачи пакета данных
	
	output wire	  load_shiftreg_o,	// Сигнал записи пакета данных в сдвиговый регистр
	output wire	  en_o,			// Выход для подтверждения валидности передаваемых последовательных данных
	output wire	  en_shiftreg_o,	// Сигнал разрешения работы сдвигового регистра
	output wire	  rst_counter_o,	// Сигнал сброса счетчика
	output wire	  busy_o,		// Сигнал занятости модуля
	output wire [7:0] data_o		// Байт данных из N-байтового буфера 
	
	);
	
	// Объявление внутренних wire/reg
	wire busy_module;	// Сигнал занятости модуля
	
	reg load_shiftreg;	// Сигнал записи пакета данных в сдвиговый регистр
	reg en_module;		// Сигнал для подтверждения валидности передаваемых последовательных данных
	reg en_shiftreg;	// Сигнал разрешения работы сдвигового регистра
	reg rst_counter;	// Сигнал сброса счетчика
	reg en_start;		// Сигнал для установки сигнала подтверждения валидности передаваемых последовательных данных
	reg en_end;		// Сигнал для сброса сигнала подтверждения валидности передаваемых последовательных данных
	reg active;		// Сигнал активности сдвигового регистра
	reg [N*8-1:0] buffer;	// N-байтовый буфер данных (FIFO)
	reg [2:0] num_byte;	// Количество байт записанных в буфер
	
	// Непрерывные присваивания  
	assign busy_module = (num_byte < N) ? 1'b0 : 1'b1; // Проверка занятости модуля
	assign load_shiftreg_o = load_shiftreg;
	assign en_o = en_module;
	assign en_shiftreg_o = en_shiftreg;
	assign rst_counter_o = rst_counter;
	assign busy_o = busy_module;
	assign data_o = buffer[7:0];
	
	always @(posedge clk_i or posedge rst_i)
	begin
		// Проверка сброса устройства
		if (rst_i)
		begin :asyn_block // Асинхронный процесс  
			buffer <= 0;		// Возвращение устройства в исходное состояние
			num_byte <= 0;
			load_shiftreg <= 1'b0;
			en_shiftreg <= 1'b0;
			en_module <= 1'b0;
			active <= 1'b0;
			en_start <= 1'b0;
			en_end <= 1'b0;
			rst_counter <= 1'b1;
		end
		else
		begin :syn_block // Синхронный процесс 
			rst_counter <= 1'b0;
			load_shiftreg <= 1'b0;
			// Проверка установки сигнала подтверждения валидности передаваемых последовательных данных
			if (en_start)
			begin
				en_module <= 1'b1;
				en_start <= 1'b0;
			end
			// Проверка сброса сигнала подтверждения валидности передаваемых последовательных данных
			if (en_end)
			begin
				en_module <= 1'b0;
				en_end <= 1'b0;
			end
			// Проверка записи в сериализатор байта данных и его занятости
			if (en_i && !busy_module)
			begin
				buffer <= buffer | (data_i << (num_byte * 8));	// Запись в буфер байта данных 
				num_byte <= num_byte + 1'b1;			// Инкремент числа байт в буфере
				// Проверка активности сдвигового регистра
				if (!active)					
				begin
					rst_counter <= 1'b1;	// Установка сигнала сброса счетчика
					load_shiftreg <= 1'b1;	// Установка сигнала загрузки пакета данных в сдвиговый регистр
					en_shiftreg <= 1'b1;	// Установка сигнала разрешения работы сдвигового регистра
					en_start <= 1'b1;	// Для установки сигнала подтверждения валидности передаваемых последовательных данных 
					active <= 1'b1;		// Установка сигнала активности сдвигового регистра
				end
			end
			// Проверка окончания передачи пакета данных
			if (count_i == 4'd11)
			begin
				buffer <= buffer >> 8;		// Сдвиг данных в буфере
				num_byte <= num_byte - 1'b1;	// Декремент числа байт в буфере
				rst_counter <= 1'b1;		// Установка сигнала сброса счетчика
				// Оценка числа байт в буфере
				if (num_byte > 3'd1)
					load_shiftreg <= 1'b1;	// Установка сигнала загрузки пакета данных в сдвиговый регистр
				else
				begin	// Если буфер опустел
					rst_counter <= 1'b1;	// Установка сигнала сброса счетчика
					en_shiftreg <= 1'b0;	// Сброс сигнала разрешения работы сдвигового регистра
					en_end <= 1'b1;		// Для сброса сигнала подтверждения валидности передаваемых последовательных данных 
					active <= 1'b0;		// Сброс сигнала активности сдвигового регистра
				end
			end
		end
	end	
	
endmodule
